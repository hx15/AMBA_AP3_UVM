`include "RTLDefines.sv"
`include "interface.sv"


package APBPackage;
   import uvm_pkg::*;

`include "uvm_macros.svh"
`include "ATransaction.sv"
`include "MSequence.sv"
`include "MSequencer.sv"
`include "MDriver.sv"
`include "MMonitor.sv"
`include "scoreboard.sv"
`include "MAgent.sv"
`include "Environment.sv"
`include "Test.sv"

endpackage // APBPackage
   
