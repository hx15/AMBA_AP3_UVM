`include "RTLDefines.sv"
`include "interface.sv"


package MPackage;
   import uvm_pkg::*;
   import common_data_types::*;
   
`include "uvm_macros.svh"
`include "MTransaction.sv"
`include "MSequence.sv"
`include "MSequencer.sv"
`include "MDriver.sv"
   
`include "MMonitor.sv"
`include "MAgent.sv"
   
endpackage // MPackage
   
   
