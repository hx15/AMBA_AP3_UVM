`include "RTLDefines.sv"
`include "interface.sv"


package EnvPackage;

   
   import uvm_pkg::*;
   import MPackage::*;
   
`include "Environment.sv"
   
`include "Test.sv"

endpackage // EnvPackage
   
   
