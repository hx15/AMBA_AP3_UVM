
package common_data_types;

typedef enum {WRTITE=0, READ=1, IDLE=2} op_type;

endpackage // data_types
   
