`include "RTLDefines.sv"
`include "interface.sv"
package APBPackage;
   import uvm_pkg::*;
   import MPackage::*;
   import EnvPackage::*;
`include "Test.sv"

endpackage // APBPackage
   
